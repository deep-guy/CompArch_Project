module DMCache(address, cache, missCount, hitCount);


endmodule